//-----------------------------------------------------------------------------
//
// Title       : Top_tb_tim
// Design      : ZegarSzachowy
// Author      : Kacper
// Company     : Tak
//
//-----------------------------------------------------------------------------
//
// File        : Top_TB_tim.v
// Generated   : Mon Jan 27 10:09:48 2025
// From        : C:\Users\Kacper\Desktop\ProjektPSC\ZegarSzachowy\src\TestBench\Top_TB_tim_settings.txt
// By          : tb_verilog.pl ver. ver 1.2s
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps
module Top_tb_tim;


//Internal signals declarations:
reg CLK;
reg CLR;
reg CE;
reg SELECT;
reg STOP;
reg Set_Impulse;
reg D1;
reg D2;
reg D3;
reg D4;
reg D5;
reg D6;
reg D7;
reg D8;
wire [6:0]seg_out;
wire [7:0]seg_select;



// Unit Under Test port map
	Top UUT (
		.CLK(CLK),
		.CLR(CLR),
		.CE(CE),
		.SELECT(SELECT),
		.STOP(STOP),
		.Set_Impulse(Set_Impulse),
		.D1(D1),
		.D2(D2),
		.D3(D3),
		.D4(D4),
		.D5(D5),
		.D6(D6),
		.D7(D7),
		.D8(D8),
		.seg_out(seg_out),
		.seg_select(seg_select));

initial
	$monitor($realtime,,"ps %h %h %h %h %h %h %h %h %h %h %h %h %h %h %h %h ",CLK,CLR,CE,SELECT,STOP,Set_Impulse,D1,D2,D3,D4,D5,D6,D7,D8,seg_out,seg_select);

//Below code was generated based on waveform file: "C:\Users\Kacper\Desktop\ProjektPSC\ZegarSzachowy\compile\Top.ver"

initial
begin : STIMUL // begin of stimulus process
	#0
	D4 = 1'b0;
	STOP = 1'b0;
	D3 = 1'b0;
	D1 = 1'b0;
	D5 = 1'b0;
	SELECT = 1'b0;
	CLR = 1'b1;
	D6 = 1'b0;
	CE = 1'b0;
	D2 = 1'b0;
	D7 = 1'b0;
	CLK = 1'b0;
	Set_Impulse = 1'b0;
	D8 = 1'b0;
    #10000; //0
	CLK = 1'b1;
    #10000; //10000
	CLK = 1'b0;
    #10000; //20000
	CLK = 1'b1;
    #10000; //30000
	CLK = 1'b0;
    #10000; //40000
	SELECT = 1'b1;
	CLR = 1'b0;
	CE = 1'b1;
	CLK = 1'b1;
    #10000; //50000
	CLK = 1'b0;
    #10000; //60000
	CLK = 1'b1;
    #10000; //70000
	CLK = 1'b0;
    #10000; //80000
	CLK = 1'b1;
    #10000; //90000
	CLK = 1'b0;
    #10000; //100000
	CLK = 1'b1;
    #10000; //110000
	CLK = 1'b0;
    #10000; //120000
	CLK = 1'b1;
    #10000; //130000
	CLK = 1'b0;
    #10000; //140000
	SELECT = 1'b0;
	CLK = 1'b1;
    #10000; //150000
	CLK = 1'b0;
    #10000; //160000
	CLK = 1'b1;
    #10000; //170000
	CLK = 1'b0;
    #10000; //180000
	CLK = 1'b1;
    #10000; //190000
	CLK = 1'b0;
    #10000; //200000
	CLK = 1'b1;
    #10000; //210000
	CLK = 1'b0;
    #10000; //220000
	CLK = 1'b1;
    #10000; //230000
	CLK = 1'b0;
    #10000; //240000
	CLK = 1'b1;
    #10000; //250000
	CLK = 1'b0;
    #10000; //260000
	CLK = 1'b1;
    #10000; //270000
	CLK = 1'b0;
    #10000; //280000
	CLK = 1'b1;
    #10000; //290000
	CLK = 1'b0;
    #10000; //300000
	CLK = 1'b1;
    #10000; //310000
	CLK = 1'b0;
    #10000; //320000
	CLK = 1'b1;
    #10000; //330000
	CLK = 1'b0;
    #10000; //340000
	SELECT = 1'b1;
	CLK = 1'b1;
    #10000; //350000
	CLK = 1'b0;
    #10000; //360000
	CLK = 1'b1;
    #10000; //370000
	CLK = 1'b0;
    #10000; //380000
	CLK = 1'b1;
    #10000; //390000
	CLK = 1'b0;
    #10000; //400000
	CLK = 1'b1;
    #10000; //410000
	CLK = 1'b0;
    #10000; //420000
	CLK = 1'b1;
    #10000; //430000
	CLK = 1'b0;
    #10000; //440000
	SELECT = 1'b0;
	CLK = 1'b1;
    #10000; //450000
	CLK = 1'b0;
    #10000; //460000
	CLK = 1'b1;
    #10000; //470000
	CLK = 1'b0;
    #10000; //480000
	CLK = 1'b1;
    #10000; //490000
	CLK = 1'b0;
    #10000; //500000
	CLK = 1'b1;
    #10000; //510000
	CLK = 1'b0;
    #10000; //520000
	CLK = 1'b1;
    #10000; //530000
	CLK = 1'b0;
    #10000; //540000
	CLK = 1'b1;
    #10000; //550000
	CLK = 1'b0;
    #10000; //560000
	CLK = 1'b1;
    #10000; //570000
	CLK = 1'b0;
    #10000; //580000
	CLK = 1'b1;
    #10000; //590000
	CLK = 1'b0;
    #10000; //600000
	CLK = 1'b1;
    #10000; //610000
	CLK = 1'b0;
    #10000; //620000
	CLK = 1'b1;
    #10000; //630000
	CLK = 1'b0;
    #10000; //640000
	CLK = 1'b1;
    #10000; //650000
	CLK = 1'b0;
    #10000; //660000
	CLK = 1'b1;
    #10000; //670000
	CLK = 1'b0;
    #10000; //680000
	CLK = 1'b1;
    #10000; //690000
	CLK = 1'b0;
    #10000; //700000
	CLK = 1'b1;
    #10000; //710000
	CLK = 1'b0;
    #10000; //720000
	CLK = 1'b1;
    #10000; //730000
	CLK = 1'b0;
    #10000; //740000
	SELECT = 1'b1;
	CLK = 1'b1;
    #10000; //750000
	CLK = 1'b0;
    #10000; //760000
	CLK = 1'b1;
    #10000; //770000
	CLK = 1'b0;
    #10000; //780000
	CLK = 1'b1;
    #10000; //790000
	SELECT = 1'b0;
	CLK = 1'b0;
    #10000; //800000
	CLK = 1'b1;
    #10000; //810000
	CLK = 1'b0;
    #10000; //820000
	CLK = 1'b1;
    #10000; //830000
	CLK = 1'b0;
    #10000; //840000
	CLK = 1'b1;
    #10000; //850000
	CLK = 1'b0;
    #10000; //860000
	CLK = 1'b1;
    #10000; //870000
	CLK = 1'b0;
    #10000; //880000
	CLK = 1'b1;
    #10000; //890000
	CLK = 1'b0;
    #10000; //900000
	CLK = 1'b1;
    #10000; //910000
	CLK = 1'b0;
    #10000; //920000
	CLK = 1'b1;
    #10000; //930000
	CLK = 1'b0;
    #10000; //940000
	STOP = 1'b1;
	SELECT = 1'b1;
	CLK = 1'b1;
    #10000; //950000
	CLK = 1'b0;
    #10000; //960000
	CLK = 1'b1;
    #10000; //970000
	CLK = 1'b0;
    #10000; //980000
	CLK = 1'b1;
    #10000; //990000
	CLK = 1'b0;
    #10000; //1000000
	CLK = 1'b1;
    #10000; //1010000
	CLK = 1'b0;
    #10000; //1020000
	CLK = 1'b1;
    #10000; //1030000
	CLK = 1'b0;
    #10000; //1040000
	D1 = 1'b1;
	CLK = 1'b1;
	Set_Impulse = 1'b1;
    #10000; //1050000
	CLK = 1'b0;
    #10000; //1060000
	D5 = 1'b1;
	CLK = 1'b1;
    #10000; //1070000
	CLK = 1'b0;
    #10000; //1080000
	D2 = 1'b1;
	CLK = 1'b1;
    #10000; //1090000
	CLK = 1'b0;
    #10000; //1100000
	D6 = 1'b1;
	CLK = 1'b1;
    #10000; //1110000
	CLK = 1'b0;
    #10000; //1120000
	D3 = 1'b1;
	CLK = 1'b1;
    #10000; //1130000
	CLK = 1'b0;
    #10000; //1140000
	D7 = 1'b1;
	CLK = 1'b1;
    #10000; //1150000
	CLK = 1'b0;
    #10000; //1160000
	D4 = 1'b1;
	CLK = 1'b1;
    #10000; //1170000
	CLK = 1'b0;
    #10000; //1180000
	CLK = 1'b1;
	D8 = 1'b1;
    #10000; //1190000
	CLK = 1'b0;
    #10000; //1200000
	CLK = 1'b1;
    #10000; //1210000
	CLK = 1'b0;
    #10000; //1220000
	CLK = 1'b1;
    #10000; //1230000
	CLK = 1'b0;
    #10000; //1240000
	CLK = 1'b1;
    #10000; //1250000
	CLK = 1'b0;
    #10000; //1260000
	CLK = 1'b1;
    #10000; //1270000
	CLK = 1'b0;
    #10000; //1280000
	CLK = 1'b1;
    #10000; //1290000
	CLK = 1'b0;
    #10000; //1300000
	CLK = 1'b1;
    #10000; //1310000
	CLK = 1'b0;
    #10000; //1320000
	CLK = 1'b1;
    #10000; //1330000
	CLK = 1'b0;
    #10000; //1340000
	STOP = 1'b0;
	D1 = 1'b0;
	CLK = 1'b1;
	Set_Impulse = 1'b0;
    #10000; //1350000
	CLK = 1'b0;
    #10000; //1360000
	CLK = 1'b1;
    #10000; //1370000
	CLK = 1'b0;
    #10000; //1380000
	CLK = 1'b1;
    #10000; //1390000
	CLK = 1'b0;
    #10000; //1400000
	CLK = 1'b1;
    #10000; //1410000
	CLK = 1'b0;
    #10000; //1420000
	CLK = 1'b1;
    #10000; //1430000
	CLK = 1'b0;
    #10000; //1440000
	CLK = 1'b1;
    #10000; //1450000
	CLK = 1'b0;
    #10000; //1460000
	CLK = 1'b1;
    #10000; //1470000
	CLK = 1'b0;
    #10000; //1480000
	CLK = 1'b1;
    #10000; //1490000
	CLK = 1'b0;
    #10000; //1500000
	CLK = 1'b1;
    #10000; //1510000
	CLK = 1'b0;
    #10000; //1520000
	CLK = 1'b1;
    #10000; //1530000
	CLK = 1'b0;
    #10000; //1540000
	CLK = 1'b1;
    #10000; //1550000
	CLK = 1'b0;
    #10000; //1560000
	CLK = 1'b1;
    #10000; //1570000
	CLK = 1'b0;
    #10000; //1580000
	CLK = 1'b1;
    #10000; //1590000
	CLK = 1'b0;
    #10000; //1600000
	CLK = 1'b1;
    #10000; //1610000
	CLK = 1'b0;
    #10000; //1620000
	CLK = 1'b1;
    #10000; //1630000
	CLK = 1'b0;
    #10000; //1640000
	CLK = 1'b1;
    #10000; //1650000
	CLK = 1'b0;
    #10000; //1660000
	CLK = 1'b1;
    #10000; //1670000
	CLK = 1'b0;
    #10000; //1680000
	CLK = 1'b1;
    #10000; //1690000
	CLK = 1'b0;
    #10000; //1700000
	CLK = 1'b1;
    #10000; //1710000
	CLK = 1'b0;
    #10000; //1720000
	CLK = 1'b1;
    #10000; //1730000
	CLK = 1'b0;
    #10000; //1740000
	CLK = 1'b1;
    #10000; //1750000
	CLK = 1'b0;
    #10000; //1760000
	CLK = 1'b1;
    #10000; //1770000
	CLK = 1'b0;
    #10000; //1780000
	CLK = 1'b1;
    #10000; //1790000
	CLK = 1'b0;
    #10000; //1800000
	CLK = 1'b1;
    #10000; //1810000
	CLK = 1'b0;
    #10000; //1820000
	CLK = 1'b1;
    #10000; //1830000
	CLK = 1'b0;
    #10000; //1840000
	CLK = 1'b1;
    #10000; //1850000
	CLK = 1'b0;
    #10000; //1860000
	CLK = 1'b1;
    #10000; //1870000
	CLK = 1'b0;
    #10000; //1880000
	CLK = 1'b1;
    #10000; //1890000
	CLK = 1'b0;
    #10000; //1900000
	CLK = 1'b1;
    #10000; //1910000
	CLK = 1'b0;
    #10000; //1920000
	CLK = 1'b1;
    #10000; //1930000
	CLK = 1'b0;
    #10000; //1940000
	CLK = 1'b1;
    #10000; //1950000
	CLK = 1'b0;
    #10000; //1960000
	CLK = 1'b1;
    #10000; //1970000
	CLK = 1'b0;
    #10000; //1980000
	CLK = 1'b1;
    #10000; //1990000
	CLK = 1'b0;
end // end of stimulus process
	



endmodule
